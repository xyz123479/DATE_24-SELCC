module SEC_DAEC_TAEC_encoder(input [63:0] message, output [71:0] codeword);

    assign codeword[71:8] = message[63:0];
    assign codeword[7] = ^(message&64'b1000000010101010000101000101010010001100000100100011010100101010);
    assign codeword[6] = ^(message&64'b0100000001010001100000100100000111011011111001010100000100010001);
    assign codeword[5] = ^(message&64'b0010000010000100010000010001110100110010000101001001001101110100);
    assign codeword[4] = ^(message&64'b0001000001001000001010001101000001000101010010100100100011100010);
    assign codeword[3] = ^(message&64'b0000100000100100100000000010010101100000101010001000100101000111);
    assign codeword[2] = ^(message&64'b0000010000010010010010000000001000101010100100110110010010010100);
    assign codeword[1] = ^(message&64'b0000001000000001001001010000000010010100010010010001011001011001);
    assign codeword[0] = ^(message&64'b0000000100000000000100101010101000000001001001001010101010111110);

endmodule