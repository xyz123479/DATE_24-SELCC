module SCC_8LC_syndrome_gen(input [71:0] codeword, output [7:0] syndrome);

    assign syndrome[7] = ^(codeword&72'b0110010111111011110011010100010111010111101101111101001000111000_10000000);
    assign syndrome[6] = ^(codeword&72'b0011001011111101111001100010001011101011110110111110100100011100_01000000);
    assign syndrome[5] = ^(codeword&72'b1001100101111110111100110001000101110101111011010111010010001110_00100000);
    assign syndrome[4] = ^(codeword&72'b1100110010111111011110010000100010111010111101100011101001000111_00010000);
    assign syndrome[3] = ^(codeword&72'b0000001110100100011100011100000110001010110011001100111100011011_00001000);
    assign syndrome[2] = ^(codeword&72'b1110010000101001111101011010010100010010110100010011010110110101_00000100);
    assign syndrome[1] = ^(codeword&72'b1001011111101111001101110001011101011110110111110100100011100010_00000010);
    assign syndrome[0] = ^(codeword&72'b1100101111110111100110111000101110101111011011111010010001110001_00000001);

endmodule
