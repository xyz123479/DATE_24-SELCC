module SEC_DED_encoder(input [63:0] message, output [71:0] codeword);

    assign codeword[71:8] = message[63:0];
    assign codeword[7] = ^(message&64'b1000101001001001001010101001001001010100101010010010100100100010);
    assign codeword[6] = ^(message&64'b0010001001001001001001010100100100101010010101001111110001001000);
    assign codeword[5] = ^(message&64'b0001001000100100100101001010100100100101001001010010001111111111);
    assign codeword[4] = ^(message&64'b0100010001000100100100100101010010100100100100101001001001001001);
    assign codeword[3] = ^(message&64'b0100100100100100010010010010011110010010100100100100100100100100);
    assign codeword[2] = ^(message&64'b0100100100100010001001001001001001001001010010100101001001111111);
    assign codeword[1] = ^(message&64'b0100100100010001000100100100100010010010010010010010010010011111);
    assign codeword[0] = ^(message&64'b0100100010001000100010010010010001001001001001001010010011100111);

endmodule