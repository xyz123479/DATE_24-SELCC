module SEC_DAEC_encoder(input [63:0] message, output [71:0] codeword);

    assign codeword[71:8] = message[63:0];
    assign codeword[7] = ^(message&64'b1001010111010110010100100100001011000100110010001101000011100000);
    assign codeword[6] = ^(message&64'b1011100110000010101001001000010110001001100100011010000111000001);
    assign codeword[5] = ^(message&64'b0110101010111010110010010000101100010011001000110100001110000011);
    assign codeword[4] = ^(message&64'b1111011001011001100100101001011000100110010001101000011000000111);
    assign codeword[3] = ^(message&64'b1001011000111101101001010010110001001100100011000000110100001110);
    assign codeword[2] = ^(message&64'b1110110011111101110010100101100010011000000110010001101000011100);
    assign codeword[1] = ^(message&64'b0110101101101111000101001011000000110001001100100011010000111000);
    assign codeword[0] = ^(message&64'b0101111011100111001010010110000101100010011001000110100001110000);

endmodule