module SCC_4LC_encoder(input [63:0] message, output [70:0] codeword);

    assign codeword[70:7] = message[63:0];
    assign codeword[6] = ^(message&64'b0001010001001100100110011110111010010110011100010111000001111101);
    assign codeword[5] = ^(message&64'b0111001110101010110101010001000111011101011010011100100001000011);
    assign codeword[4] = ^(message&64'b0011000010011011111100110110011001111000111001011001010001011100);
    assign codeword[3] = ^(message&64'b1000111000101111111110011011001100111100010100101100101000101110);
    assign codeword[2] = ^(message&64'b1100110011110101111111001101100110011110001010010110010100010111);
    assign codeword[1] = ^(message&64'b0000101001110110011001111000101001011001010001011100001011110110);
    assign codeword[0] = ^(message&64'b0101010100011001001100111100110100101100101000101110000111111011);

endmodule