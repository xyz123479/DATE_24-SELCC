module SCC_8LC_encoder(input [63:0] message, output [71:0] codeword);

    assign codeword[71:8] = message[63:0];
    assign codeword[7] = ^(message&64'b0110010111111011110011010100010111010111101101111101001000111000);
    assign codeword[6] = ^(message&64'b0011001011111101111001100010001011101011110110111110100100011100);
    assign codeword[5] = ^(message&64'b1001100101111110111100110001000101110101111011010111010010001110);
    assign codeword[4] = ^(message&64'b1100110010111111011110010000100010111010111101100011101001000111);
    assign codeword[3] = ^(message&64'b0000001110100100011100011100000110001010110011001100111100011011);
    assign codeword[2] = ^(message&64'b1110010000101001111101011010010100010010110100010011010110110101);
    assign codeword[1] = ^(message&64'b1001011111101111001101110001011101011110110111110100100011100010);
    assign codeword[0] = ^(message&64'b1100101111110111100110111000101110101111011011111010010001110001);

endmodule